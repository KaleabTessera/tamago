module tamago.aca.bank;


service Deposit {

	refine service ACASecurity in tamago.aca.core;
	
	method void init() {
		id init;
	}
	
	method void deposit(int clid, int cid,tamago.ext.aca2.ACA aca) {
	       id deposit;
	}
	method void cancel(int clid, int cid,tamago.ext.aca2.ACA aca) {
	       id cancel;
	}
	method void validate(int clid, int cid,tamago.ext.aca2.ACA aca) {
		id validate;
	}
	method void validate_director(int clid, int cid,tamago.ext.aca2.ACA aca) {
		id validate_dir;
	}
	
	method void check(int clid, int cid,tamago.ext.aca2.ACA aca) {
		id check;
		//verifie que le client est ok
		// cheque en bois
	}
	
	method void register(int clid, int cid,tamago.ext.aca2.ACA aca) {
		id register;
		// historique de la banque
	}
}
