module tamago.aca.bank;

service Cheque {

}