module tamago.aca.bank;

service DepositService {
	refine service ACASecurity in tamago.aca.core;
	property read int opNumber;
	
	method void init() {
		id init;
		post (#opNumber < 0);
	}
	
	method void deposit(tamago.ext.aca2.ACA aca) {
		id deposit;
	}
	method void cancel(tamago.ext.aca2.ACA aca) {
		id cancel;
	}
	method void validate(tamago.ext.aca2.ACA aca) {
		id validate;
	}
	method void validate_director(tamago.ext.aca2.ACA aca) {
		id validate_dir;
	}
	method void check(tamago.ext.aca2.ACA aca) {
		id check;
		post (#opNumber > 0);
	}

	method void register(tamago.ext.aca2.ACA aca) {
		id register;
		post (#opNumber > 0);
	}
	
	behavior {
		default state ninit;
		states {
			state ninit {
				allow init;
			}
			state initialized {
				allow deposit;
			}
			state deposed {
				allow check;
				allow register;
			}
			state checked {
				allow register;
			}
			state registered {
				allow check;
			}
			state waited {
				allow validate;
				allow validate_dir;
				allow cancel;
			}
			state validated {
				allow validate_dir;
			}
			state validateDir {
				allow validate;
			}
			state cancelled {
				allow init;
			}
			state completed {
				allow init;
			}
		}
		transitions {
			transition from ninit to initialized with init;
			transition from initialized to deposed with deposit;
			transition from deposed to checked with check;
			transition from deposed to registered with register;
			transition from checked to waited with register;
			transition from registered to waited with check;
			transition from waited to validated with validate;
			transition from waited to validateDir with validate_dir;
			transition from waited to cancelled with cancel;
			transition from validated to completed with validate_dir;
			transition from validateDir to completed with validate;
			transition from cancelled to initialized with init;
			transition from completed to initialized with init;
		}
	}
	
}