module tamago.aca.bank;


service Bank {
}