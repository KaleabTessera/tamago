module tamago.aca;

component VBanqueComp {
    provide service VBanque in tamago.aca;
}
