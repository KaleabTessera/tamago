module tamago.aca.core;


service ACASecurity {
	property readwrite bool acaInitialised;
	
	method void init() {
		id acasecurity_init;
		post acaInitialised;
	}
}