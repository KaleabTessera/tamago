module org.tamago.example;



component CompBucket {
	provide service Bucket in org.tamago.example;
		
	require service Bucket in org.tamago.example as a;
	require service Bucket in org.tamago.example as b;
	require service Bucket in org.tamago.example as c;
		
	method void foo() {
		id qqchose;
		//pre ((3+2) > 1);
	}
	
}