module tamago.aca.bank;


service Client {

}