module org.tamago.example;

using java.lang.*;

service Bucket {
	property read int quantity;
	method void foo(int a) {
        id foo;
		//post 4+3 == 7;
	}
	
	behavior {
		default state toto;
		states {
			state toto { allow foo; }
		}
		transitions {
			transition from toto to toto with foo when true;
		}
	}
}