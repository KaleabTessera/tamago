module org.tamago.example;

using java.lang.String;

service Bucket {
	property read int quantity;
	method void foo(int a) {
		id foo;
		//pre @instate(toto);
	}
	
	behavior {
		default state toto;
		states {
			state toto { allow foo; }
		}
		transitions {
			transition from toto to toto with foo when true;
		}
	}
}