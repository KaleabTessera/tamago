module tamago.aca.bank;


service Deposit {
	
	method void deposit(int clid, int cid,tamago.ext.aca2.ACA aca) {
	       id deposit;
	}
	method void cancel(int clid, int cid,tamago.ext.aca2.ACA aca) {
	       id cancel;
	}
	method void validate(int clid, int cid,tamago.ext.aca2.ACA aca) {
		id validate;
	}
	method void validate_director(int clid, int cid,tamago.ext.aca2.ACA aca) {
		id validate_dir;
	}
	
	method void check(int clid, int cid,tamago.ext.aca2.ACA aca) {
		id check;
	}
	
	method void register(int clid, int cid,tamago.ext.aca2.ACA aca) {
		id register;
	}
}
