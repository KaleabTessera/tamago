module tamago.aca.bank;


service Deposit {

	refine service ACASecurity in tamago.aca.core;
	
	property read int opNumber; // numero d'ordre
	
	
	method void init() {
		id init;
	}
	
	method void deposit(tamago.ext.aca2.ACA aca) {
	       id deposit;
	}
	method void cancel(tamago.ext.aca2.ACA aca) {
	       id cancel;
	}
	method void validate(tamago.ext.aca2.ACA aca) {
		id validate;
	}
	method void validate_director(tamago.ext.aca2.ACA aca) {
		id validate_dir;
	}
	
	method void check(tamago.ext.aca2.ACA aca) {
		id check;
		//verifie que le client est ok
		// cheque en bois
	}
	
	method void register(tamago.ext.aca2.ACA aca) {
		id register;
		// historique de la banque
	}
	
	behavior {
		default state ninit;
		states {
		state ninit {
			allow init;
		}
		state initialized {
			allow deposit;
		}
		state deposed {
			allow check;
			allow register;
		}
		state checked {
			allow register;
		}
		state registered {
			allow check;
		}
		state checkedregistered {
			allow cancel;
			allow validate;
			allow validate_dir;
		}
		
		state cancelled {
			allow init;
		}
		state validated {
			allow validate_dir;
		}
		state validatedDir {
			allow validate;
		}
		}
		transitions {
			transition from ninit to initialized with init;
			transition from initialized to deposed with deposit;
			transition from deposed to checked with check;
			transition from deposed to registered with register;
			transition from checked to checkedregistered with register;
			transition from registered to checkedregistered with check;
			transition from checkedregistered to cancelled with cancel;
			transition from checkedregistered to validated with validate;
			transition from checkedregistered to validatedDir with validate_dir;
		}
	}
}
